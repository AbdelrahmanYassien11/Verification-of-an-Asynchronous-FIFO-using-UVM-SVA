class env_config;
	virtual inf env_config_my_vif;

	function new(virtual inf env_config_my_vif);
    	this.env_config_my_vif = env_config_my_vif;
 	endfunction : new
endclass : env_config

