interface inf(input clk);


logic rst_n, d;
logic q;


endinterface : inf